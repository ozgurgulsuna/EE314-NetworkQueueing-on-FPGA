module buffer(
	input clk,
	input [3:0] sw_in,
);