library verilog;
use verilog.vl_types.all;
entity buffer_vlg_vec_tst is
end buffer_vlg_vec_tst;
