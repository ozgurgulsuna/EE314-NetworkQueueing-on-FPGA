library verilog;
use verilog.vl_types.all;
entity decision_test_vlg_vec_tst is
end decision_test_vlg_vec_tst;
