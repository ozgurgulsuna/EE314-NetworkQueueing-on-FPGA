library verilog;
use verilog.vl_types.all;
entity switch_sim_vlg_vec_tst is
end switch_sim_vlg_vec_tst;
