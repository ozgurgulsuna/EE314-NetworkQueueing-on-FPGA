library verilog;
use verilog.vl_types.all;
entity clk_div_vlg_vec_tst is
end clk_div_vlg_vec_tst;
