library verilog;
use verilog.vl_types.all;
entity debouncer_vlg_vec_tst is
end debouncer_vlg_vec_tst;
