library verilog;
use verilog.vl_types.all;
entity button_test_vlg_vec_tst is
end button_test_vlg_vec_tst;
