library verilog;
use verilog.vl_types.all;
entity buffer_sim_vlg_vec_tst is
end buffer_sim_vlg_vec_tst;
